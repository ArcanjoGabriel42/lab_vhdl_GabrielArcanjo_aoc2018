library ieee;
use ieee.std_logic_1164.all;

Entity Mux_4 is
	Port
	(
		A,B,C,D: in std_logic_vector(15 downto 0);
		Output: out std_logic_vector(15 downto 0);
		Se: in std_logic_vector(1 downto 0)
	);
End Mux_4;

Architecture behavior of Mux_4 is 
Begin
	Process(A,B,C,D,Se)
	Begin
		Case Se is
			when "00" => Output <= A;
			when "01" => Output <= B;
			when "10" => Output <= C;
			when "11" => Output <= D;

			when others => Output <= "ZZZZZZZZZZZZZZZZ";
		End Case;
	End Process;
End behavior;